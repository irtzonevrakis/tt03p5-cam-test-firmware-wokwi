// A simple associative array in verilog: Main array logic.
// Copyright (C) 2023 Ioannis-Rafail Tzonevrakis.


module wokwi(input wire ui_in_0,
             input wire ui_in_1,
             input wire ui_in_2,
             input wire ui_in_3,
             input wire ui_in_4,
             input wire ui_in_5,
             input wire ui_in_6,
             input wire ui_in_7,
             output wire uo_out_0,
             output wire uo_out_1,
             output wire uo_out_2,
             output wire uo_out_3,
             output wire uo_out_4,
             output wire uo_out_5,
             output wire uo_out_6,
             output wire uo_out_7,
	     output wire uio_in_0,
	     output wire uio_in_1,
	     output wire uio_in_2,
	     output wire uio_in_3,
	     output wire uio_in_4,
	     output wire uio_in_5,
	     output wire uio_in_6,
	     output wire uio_in_7,
             output wire uio_out_0,
             output wire uio_out_1,
             output wire uio_out_2,
             output wire uio_out_3,
             output wire uio_out_4,
             output wire uio_out_5,
             output wire uio_out_6,
             output wire uio_out_7,
             input  wire ena,
             input  wire clk,
             input  wire rst_n);
  
  wire [7:0] uio_oe;
  
  tt_um_cam cam0 (.clk(clk), 
                  .ena(ena), 
                  .rst_n(rst_n),
                  .ui_in({ui_in_7,
                          ui_in_6,
                          ui_in_5,
                          ui_in_4,
                          ui_in_3,
                          ui_in_2,
                          ui_in_1,
                          ui_in_0}),
                  .uo_out({uo_out_7,
                           uo_out_6,
                           uo_out_5,
                           uo_out_4,
                           uo_out_3,
                           uo_out_2,
                           uo_out_1,
                           uo_out_0}),
                  .uio_in({uio_in_7,
                           uio_in_6,
                           uio_in_5,
                           uio_in_4,
                           uio_in_3,
                           uio_in_2,
                           uio_in_1,
                           uio_in_0}),
                 .uio_out({uio_out_7,
                           uio_out_6,
                           uio_out_5,
                           uio_out_4,
                           uio_out_3,
                           uio_out_2,
                           uio_out_1,
                           uio_out_0}),
                 .uio_oe(uio_oe));
endmodule
